module xdma_gen3_x1_minimal (
    input PCIE_REFCLK1_N,
    input PCIE_REFCLK1_P,
    input SYSCLK2_N,
    input SYSCLK2_P,
    input SYSCLK3_N,
    input SYSCLK3_P
);

endmodule
